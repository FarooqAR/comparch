module pipelined_processor (
	input clk,    // Clock
	input rst,  // Asynchronous reset active low
);
	//IF/ID

	//ID/EX

	//EX/MEM

	//MEM/WB
	
endmodule